module controller #(parameter W=32) 
    (   
        input clk,
        input [3:0] Cond,
        input [1:0] Op,
        input [5:0] Func,
        input [3:0] Rd,
        output PCSrc,
        output RegWrite,
        output MemWrite,
        output MemToReg,
        output AluSrc,
        output [1:0] ImmSrc,
        output [1:0] RegSrc,
        output [1:0] AluControl
    );




    








endmodule
